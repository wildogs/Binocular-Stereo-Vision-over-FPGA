
wire kernel_monitor_reset;
wire kernel_monitor_clock;
wire kernel_monitor_report;
assign kernel_monitor_reset = ~ap_rst_n;
assign kernel_monitor_clock = ap_clk;
assign kernel_monitor_report = 1'b0;
wire [6:0] axis_block_sigs;
wire [40:0] inst_idle_sigs;
wire [29:0] inst_block_sigs;
wire kernel_block;

assign axis_block_sigs[0] = ~AXIvideo2xfMat_8_0_600_800_1_2_1_U0.grp_AXIvideo2xfMat_8_0_600_800_1_2_1_Pipeline_loop_start_hunt_fu_185.vid_inL_TDATA_blk_n;
assign axis_block_sigs[1] = ~AXIvideo2xfMat_8_0_600_800_1_2_1_U0.grp_AXIvideo2xfMat_8_0_600_800_1_2_1_Pipeline_loop_col_zxi2mat_fu_205.vid_inL_TDATA_blk_n;
assign axis_block_sigs[2] = ~AXIvideo2xfMat_8_0_600_800_1_2_1_U0.grp_AXIvideo2xfMat_8_0_600_800_1_2_1_Pipeline_loop_last_hunt_fu_232.vid_inL_TDATA_blk_n;
assign axis_block_sigs[3] = ~AXIvideo2xfMat_8_0_600_800_1_2_U0.grp_AXIvideo2xfMat_8_0_600_800_1_2_Pipeline_loop_start_hunt_fu_185.vid_inR_TDATA_blk_n;
assign axis_block_sigs[4] = ~AXIvideo2xfMat_8_0_600_800_1_2_U0.grp_AXIvideo2xfMat_8_0_600_800_1_2_Pipeline_loop_col_zxi2mat_fu_205.vid_inR_TDATA_blk_n;
assign axis_block_sigs[5] = ~AXIvideo2xfMat_8_0_600_800_1_2_U0.grp_AXIvideo2xfMat_8_0_600_800_1_2_Pipeline_loop_last_hunt_fu_232.vid_inR_TDATA_blk_n;
assign axis_block_sigs[6] = ~xfMat2AXIvideo_8_0_600_800_1_2_U0.grp_xfMat2AXIvideo_8_0_600_800_1_2_Pipeline_loop_col_mat2axi_fu_86.vid_out_TDATA_blk_n;

assign inst_idle_sigs[0] = Loop_VITIS_LOOP_46_1_proc_U0.ap_idle;
assign inst_block_sigs[0] = (Loop_VITIS_LOOP_46_1_proc_U0.ap_done & ~Loop_VITIS_LOOP_46_1_proc_U0.ap_continue);
assign inst_idle_sigs[1] = Loop_VITIS_LOOP_55_2_proc_U0.ap_idle;
assign inst_block_sigs[1] = (Loop_VITIS_LOOP_55_2_proc_U0.ap_done & ~Loop_VITIS_LOOP_55_2_proc_U0.ap_continue);
assign inst_idle_sigs[2] = Block_for_end72_proc_U0.ap_idle;
assign inst_block_sigs[2] = (Block_for_end72_proc_U0.ap_done & ~Block_for_end72_proc_U0.ap_continue);
assign inst_idle_sigs[3] = AXIvideo2xfMat_8_0_600_800_1_2_1_U0.ap_idle;
assign inst_block_sigs[3] = (AXIvideo2xfMat_8_0_600_800_1_2_1_U0.ap_done & ~AXIvideo2xfMat_8_0_600_800_1_2_1_U0.ap_continue) | ~AXIvideo2xfMat_8_0_600_800_1_2_1_U0.grp_AXIvideo2xfMat_8_0_600_800_1_2_1_Pipeline_loop_col_zxi2mat_fu_205.imgL_in_data_blk_n | ~AXIvideo2xfMat_8_0_600_800_1_2_1_U0.imgL_in_rows_c_blk_n | ~AXIvideo2xfMat_8_0_600_800_1_2_1_U0.imgL_in_cols_c_blk_n;
assign inst_idle_sigs[4] = AXIvideo2xfMat_8_0_600_800_1_2_U0.ap_idle;
assign inst_block_sigs[4] = (AXIvideo2xfMat_8_0_600_800_1_2_U0.ap_done & ~AXIvideo2xfMat_8_0_600_800_1_2_U0.ap_continue) | ~AXIvideo2xfMat_8_0_600_800_1_2_U0.grp_AXIvideo2xfMat_8_0_600_800_1_2_Pipeline_loop_col_zxi2mat_fu_205.imgR_in_data_blk_n | ~AXIvideo2xfMat_8_0_600_800_1_2_U0.imgR_in_rows_c_blk_n | ~AXIvideo2xfMat_8_0_600_800_1_2_U0.imgR_in_cols_c_blk_n;
assign inst_idle_sigs[5] = InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0.ap_idle;
assign inst_block_sigs[5] = (InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0.ap_done & ~InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0.ap_continue) | ~InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0.grp_xFInitUndistortRectifyMapInverseKernel_fu_40.grp_xFInitUndistortRectifyMapInverseKernel_Pipeline_loop_height_loop_width_fu_152.mapxRMat_data_blk_n | ~InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0.grp_xFInitUndistortRectifyMapInverseKernel_fu_40.grp_xFInitUndistortRectifyMapInverseKernel_Pipeline_loop_height_loop_width_fu_152.mapyRMat_data_blk_n;
assign inst_idle_sigs[6] = remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.ap_idle;
assign inst_block_sigs[6] = (remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.ap_done & ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.ap_continue) | ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_Block_entry1_proc_U0.p_src_mat_rows_blk_n | ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_Block_entry1_proc_U0.p_src_mat_cols_blk_n | ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_Pipeline_loop_width_fu_104.imgL_in_data_blk_n | ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_Pipeline_loop_width_fu_104.leftRemappedMat_data_blk_n | ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_Pipeline_loop_width_fu_104.mapxLMat_data_blk_n | ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_Pipeline_loop_width_fu_104.mapyLMat_data_blk_n;
assign inst_idle_sigs[7] = InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0.ap_idle;
assign inst_block_sigs[7] = (InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0.ap_done & ~InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0.ap_continue) | ~InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0.grp_xFInitUndistortRectifyMapInverseKernel_fu_40.grp_xFInitUndistortRectifyMapInverseKernel_Pipeline_loop_height_loop_width_fu_152.mapxRMat_data_blk_n | ~InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0.grp_xFInitUndistortRectifyMapInverseKernel_fu_40.grp_xFInitUndistortRectifyMapInverseKernel_Pipeline_loop_height_loop_width_fu_152.mapyRMat_data_blk_n;
assign inst_idle_sigs[8] = remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.ap_idle;
assign inst_block_sigs[8] = (remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.ap_done & ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.ap_continue) | ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_Block_entry1_proc_U0.p_src_mat_rows_blk_n | ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_Block_entry1_proc_U0.p_src_mat_cols_blk_n | ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_Pipeline_loop_width_fu_104.imgR_in_data_blk_n | ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_Pipeline_loop_width_fu_104.rightRemappedMat_data_blk_n | ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_Pipeline_loop_width_fu_104.mapxRMat_data_blk_n | ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_Pipeline_loop_width_fu_104.mapyRMat_data_blk_n;
assign inst_idle_sigs[9] = StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.ap_idle;
assign inst_block_sigs[9] = (StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.ap_done & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.ap_continue) | ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0.grp_xFSobelFilter3x3_0_3_600_800_1_0_4_1_2_2_2_1_6_800_false_s_fu_36.grp_xFSobelFilter3x3_Pipeline_Clear_Row_Loop_fu_148.rightRemappedMat_data_blk_n | ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0.grp_xFSobelFilter3x3_0_3_600_800_1_0_4_1_2_2_2_1_6_800_false_s_fu_36.grp_xFSobelFilter3x3_Pipeline_Col_Loop_fu_157.rightRemappedMat_data_blk_n | ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_U0.grp_xFSobelFilter3x3_0_3_600_800_1_0_4_1_2_2_2_1_6_800_false_s_fu_36.grp_xFSobelFilter3x3_Pipeline_Clear_Row_Loop_fu_148.rightRemappedMat_data_blk_n | ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_U0.grp_xFSobelFilter3x3_0_3_600_800_1_0_4_1_2_2_2_1_6_800_false_s_fu_36.grp_xFSobelFilter3x3_Pipeline_Col_Loop_fu_157.rightRemappedMat_data_blk_n | ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0.grp_xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_Pipeline_VITIS_LOOP_fu_46.img_disp16u_data_blk_n;
assign inst_idle_sigs[10] = Block_for_end7235_proc_U0.ap_idle;
assign inst_block_sigs[10] = (Block_for_end7235_proc_U0.ap_done & ~Block_for_end7235_proc_U0.ap_continue);
assign inst_idle_sigs[11] = ConvertShiftAbs_U0.ap_idle;
assign inst_block_sigs[11] = (ConvertShiftAbs_U0.ap_done & ~ConvertShiftAbs_U0.ap_continue) | ~ConvertShiftAbs_U0.grp_ConvertShiftAbs_Pipeline_loop_width_fu_38.img_disp16u_data_blk_n | ~ConvertShiftAbs_U0.grp_ConvertShiftAbs_Pipeline_loop_width_fu_38.img_disp8u_data_blk_n;
assign inst_idle_sigs[12] = Block_for_end7237_proc_U0.ap_idle;
assign inst_block_sigs[12] = (Block_for_end7237_proc_U0.ap_done & ~Block_for_end7237_proc_U0.ap_continue);
assign inst_idle_sigs[13] = erode_0_0_600_800_0_3_3_1_1_2_2_U0.ap_idle;
assign inst_block_sigs[13] = (erode_0_0_600_800_0_3_3_1_1_2_2_U0.ap_done & ~erode_0_0_600_800_0_3_3_1_1_2_2_U0.ap_continue) | ~erode_0_0_600_800_0_3_3_1_1_2_2_U0.grp_xferode_600_800_1_0_1_2_2_0_801_3_3_s_fu_34.grp_xferode_600_800_1_0_1_2_2_0_801_3_3_Pipeline_Col_Loop_fu_155.img_disp8u_data_blk_n | ~erode_0_0_600_800_0_3_3_1_1_2_2_U0.grp_xferode_600_800_1_0_1_2_2_0_801_3_3_s_fu_34.grp_xferode_600_800_1_0_1_2_2_0_801_3_3_Pipeline_VITIS_LOOP_298_2_fu_146.img_disp8u_data_blk_n | ~erode_0_0_600_800_0_3_3_1_1_2_2_U0.grp_xferode_600_800_1_0_1_2_2_0_801_3_3_s_fu_34.grp_xferode_600_800_1_0_1_2_2_0_801_3_3_Pipeline_Col_Loop_fu_155.img_disp8u_erode_data_blk_n;
assign inst_idle_sigs[14] = Block_for_end7239_proc_U0.ap_idle;
assign inst_block_sigs[14] = (Block_for_end7239_proc_U0.ap_done & ~Block_for_end7239_proc_U0.ap_continue);
assign inst_idle_sigs[15] = dilate_0_0_600_800_0_3_3_1_1_2_2_U0.ap_idle;
assign inst_block_sigs[15] = (dilate_0_0_600_800_0_3_3_1_1_2_2_U0.ap_done & ~dilate_0_0_600_800_0_3_3_1_1_2_2_U0.ap_continue) | ~dilate_0_0_600_800_0_3_3_1_1_2_2_U0.grp_xfdilate_600_800_1_0_1_2_2_0_801_3_3_s_fu_34.grp_xfdilate_600_800_1_0_1_2_2_0_801_3_3_Pipeline_Col_Loop_fu_155.img_disp8u_erode_data_blk_n | ~dilate_0_0_600_800_0_3_3_1_1_2_2_U0.grp_xfdilate_600_800_1_0_1_2_2_0_801_3_3_s_fu_34.grp_xfdilate_600_800_1_0_1_2_2_0_801_3_3_Pipeline_VITIS_LOOP_294_2_fu_146.img_disp8u_erode_data_blk_n | ~dilate_0_0_600_800_0_3_3_1_1_2_2_U0.grp_xfdilate_600_800_1_0_1_2_2_0_801_3_3_s_fu_34.grp_xfdilate_600_800_1_0_1_2_2_0_801_3_3_Pipeline_Col_Loop_fu_155.img_disp8u_dilate_data_blk_n;
assign inst_idle_sigs[16] = xfMat2AXIvideo_8_0_600_800_1_2_U0.ap_idle;
assign inst_block_sigs[16] = (xfMat2AXIvideo_8_0_600_800_1_2_U0.ap_done & ~xfMat2AXIvideo_8_0_600_800_1_2_U0.ap_continue) | ~xfMat2AXIvideo_8_0_600_800_1_2_U0.grp_xfMat2AXIvideo_8_0_600_800_1_2_Pipeline_loop_col_mat2axi_fu_86.img_disp8u_dilate_data_blk_n;
assign inst_idle_sigs[17] = remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_Block_entry1_proc_U0.ap_idle;
assign inst_block_sigs[17] = (remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_Block_entry1_proc_U0.ap_done & ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_Block_entry1_proc_U0.ap_continue);
assign inst_idle_sigs[18] = remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0.ap_idle;
assign inst_block_sigs[18] = (remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0.ap_done & ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0.ap_continue);
assign inst_idle_sigs[19] = remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_Block_entry1_proc_U0.ap_idle;
assign inst_block_sigs[19] = (remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_Block_entry1_proc_U0.ap_done & ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_Block_entry1_proc_U0.ap_continue);
assign inst_idle_sigs[20] = remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0.ap_idle;
assign inst_block_sigs[20] = (remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0.ap_done & ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0.ap_continue);
assign inst_idle_sigs[21] = StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.ap_idle;
assign inst_block_sigs[21] = (StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.ap_done & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.ap_continue);
assign inst_idle_sigs[22] = StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0.ap_idle;
assign inst_block_sigs[22] = (StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0.ap_done & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0.ap_continue);
assign inst_idle_sigs[23] = StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0.ap_idle;
assign inst_block_sigs[23] = (StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0.ap_done & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0.ap_continue);
assign inst_idle_sigs[24] = StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0.ap_idle;
assign inst_block_sigs[24] = (StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0.ap_done & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0.ap_continue);
assign inst_idle_sigs[25] = StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_U0.ap_idle;
assign inst_block_sigs[25] = (StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_U0.ap_done & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_U0.ap_continue);
assign inst_idle_sigs[26] = StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0.ap_idle;
assign inst_block_sigs[26] = (StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0.ap_done & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0.ap_continue);
assign inst_idle_sigs[27] = StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0.ap_idle;
assign inst_block_sigs[27] = (StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0.ap_done & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0.ap_continue);
assign inst_idle_sigs[28] = StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0.ap_idle;
assign inst_block_sigs[28] = (StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0.ap_done & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0.ap_continue);
assign inst_idle_sigs[29] = StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0.ap_idle;
assign inst_block_sigs[29] = (StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0.ap_done & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0.ap_continue);

assign inst_idle_sigs[30] = 1'b0;
assign inst_idle_sigs[31] = AXIvideo2xfMat_8_0_600_800_1_2_1_U0.ap_idle;
assign inst_idle_sigs[32] = AXIvideo2xfMat_8_0_600_800_1_2_1_U0.grp_AXIvideo2xfMat_8_0_600_800_1_2_1_Pipeline_loop_start_hunt_fu_185.ap_idle;
assign inst_idle_sigs[33] = AXIvideo2xfMat_8_0_600_800_1_2_1_U0.grp_AXIvideo2xfMat_8_0_600_800_1_2_1_Pipeline_loop_col_zxi2mat_fu_205.ap_idle;
assign inst_idle_sigs[34] = AXIvideo2xfMat_8_0_600_800_1_2_1_U0.grp_AXIvideo2xfMat_8_0_600_800_1_2_1_Pipeline_loop_last_hunt_fu_232.ap_idle;
assign inst_idle_sigs[35] = AXIvideo2xfMat_8_0_600_800_1_2_U0.ap_idle;
assign inst_idle_sigs[36] = AXIvideo2xfMat_8_0_600_800_1_2_U0.grp_AXIvideo2xfMat_8_0_600_800_1_2_Pipeline_loop_start_hunt_fu_185.ap_idle;
assign inst_idle_sigs[37] = AXIvideo2xfMat_8_0_600_800_1_2_U0.grp_AXIvideo2xfMat_8_0_600_800_1_2_Pipeline_loop_col_zxi2mat_fu_205.ap_idle;
assign inst_idle_sigs[38] = AXIvideo2xfMat_8_0_600_800_1_2_U0.grp_AXIvideo2xfMat_8_0_600_800_1_2_Pipeline_loop_last_hunt_fu_232.ap_idle;
assign inst_idle_sigs[39] = xfMat2AXIvideo_8_0_600_800_1_2_U0.ap_idle;
assign inst_idle_sigs[40] = xfMat2AXIvideo_8_0_600_800_1_2_U0.grp_xfMat2AXIvideo_8_0_600_800_1_2_Pipeline_loop_col_mat2axi_fu_86.ap_idle;

stereolbm_axis_cambm_hls_deadlock_idx0_monitor stereolbm_axis_cambm_hls_deadlock_idx0_monitor_U (
    .clock(kernel_monitor_clock),
    .reset(kernel_monitor_reset),
    .axis_block_sigs(axis_block_sigs),
    .inst_idle_sigs(inst_idle_sigs),
    .inst_block_sigs(inst_block_sigs),
    .block(kernel_block)
);


always @ (kernel_block or kernel_monitor_reset) begin
    if (kernel_block == 1'b1 && kernel_monitor_reset == 1'b0) begin
        find_kernel_block = 1'b1;
    end
    else begin
        find_kernel_block = 1'b0;
    end
end
