   
    parameter PROC_NUM = 30;
    parameter ST_IDLE = 3'b000;
    parameter ST_FILTER_FAKE = 3'b001;
    parameter ST_DL_DETECTED = 3'b010;
    parameter ST_DL_REPORT = 3'b100;
   

    reg [2:0] CS_fsm;
    reg [2:0] NS_fsm;
    reg [PROC_NUM - 1:0] dl_detect_reg;
    reg [PROC_NUM - 1:0] dl_done_reg;
    reg [PROC_NUM - 1:0] origin_reg;
    reg [PROC_NUM - 1:0] dl_in_vec_reg;
    reg [31:0] dl_keep_cnt;
    integer i;
    integer fp;

    // FSM State machine
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            CS_fsm <= ST_IDLE;
        end
        else begin
            CS_fsm <= NS_fsm;
        end
    end
    always @ (CS_fsm or dl_in_vec or dl_detect_reg or dl_done_reg or dl_in_vec or origin_reg or dl_keep_cnt) begin
        case (CS_fsm)
            ST_IDLE : begin
                if (|dl_in_vec) begin
                    NS_fsm = ST_FILTER_FAKE;
                end
                else begin
                    NS_fsm = ST_IDLE;
                end
            end
            ST_FILTER_FAKE: begin
                if (dl_keep_cnt >= 32'd1000) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                else if (dl_detect_reg != (dl_detect_reg & dl_in_vec)) begin
                    NS_fsm = ST_IDLE;
                end
                else begin
                    NS_fsm = ST_FILTER_FAKE;
                end
            end
            ST_DL_DETECTED: begin
                // has unreported deadlock cycle
                if (dl_detect_reg != dl_done_reg) begin
                    NS_fsm = ST_DL_REPORT;
                end
                else begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
            ST_DL_REPORT: begin
                if (|(dl_in_vec & origin_reg)) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                else begin
                    NS_fsm = ST_DL_REPORT;
                end
            end
            default: NS_fsm = ST_IDLE;
        endcase
    end

    // dl_detect_reg record the procs that first detect deadlock
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_detect_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_IDLE) begin
                dl_detect_reg <= dl_in_vec;
            end
        end
    end

    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_keep_cnt <= 32'h0;
        end
        else begin
            if (CS_fsm == ST_FILTER_FAKE && (dl_detect_reg == (dl_detect_reg & dl_in_vec))) begin
                dl_keep_cnt <= dl_keep_cnt + 32'h1;
            end
            else if (CS_fsm == ST_FILTER_FAKE && (dl_detect_reg != (dl_detect_reg & dl_in_vec))) begin
                dl_keep_cnt <= 32'h0;
            end
        end
    end

    // dl_detect_out keeps in high after deadlock detected
    assign dl_detect_out = (|dl_detect_reg) && (CS_fsm == ST_DL_DETECTED || CS_fsm == ST_DL_REPORT);

    // dl_done_reg record the cycles has been reported
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_done_reg <= 'b0;
        end
        else begin
            if ((CS_fsm == ST_DL_REPORT) && (|(dl_in_vec & dl_detect_reg) == 'b1)) begin
                dl_done_reg <= dl_done_reg | dl_in_vec;
            end
        end
    end

    // clear token once a cycle is done
    assign token_clear = (CS_fsm == ST_DL_REPORT) ? ((|(dl_in_vec & origin_reg)) ? 'b1 : 'b0) : 'b0;

    // origin_reg record the current cycle start id
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            origin_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                origin_reg <= origin;
            end
        end
    end
   
    // origin will be valid for only one cycle
    wire [PROC_NUM*PROC_NUM - 1:0] origin_tmp;
    assign origin_tmp[PROC_NUM - 1:0] = (dl_detect_reg[0] & ~dl_done_reg[0]) ? 'b1 : 'b0;
    genvar j;
    generate
    for(j = 1;j < PROC_NUM;j = j + 1) begin: F1
        assign origin_tmp[j*PROC_NUM +: PROC_NUM] = (dl_detect_reg[j] & ~dl_done_reg[j]) ? ('b1 << j) : origin_tmp[(j - 1)*PROC_NUM +: PROC_NUM];
    end
    endgenerate
    always @ (CS_fsm or origin_tmp) begin
        if (CS_fsm == ST_DL_DETECTED) begin
            origin = origin_tmp[(PROC_NUM - 1)*PROC_NUM +: PROC_NUM];
        end
        else begin
            origin = 'b0;
        end
    end

    
    // dl_in_vec_reg record the current cycle dl_in_vec
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_in_vec_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                dl_in_vec_reg <= origin;
            end
            else if (CS_fsm == ST_DL_REPORT) begin
                dl_in_vec_reg <= dl_in_vec;
            end
        end
    end
    
    // find_df_deadlock to report the deadlock
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            find_df_deadlock <= 1'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED && dl_detect_reg == dl_done_reg) begin
                find_df_deadlock <= 1'b1;
            end
            else if (CS_fsm == ST_IDLE) begin
                find_df_deadlock <= 1'b0;
            end
        end
    end
    
    // get the first valid proc index in dl vector
    function integer proc_index(input [PROC_NUM - 1:0] dl_vec);
        begin
            proc_index = 0;
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_vec[i]) begin
                    proc_index = i;
                end
            end
        end
    endfunction

    // get the proc path based on dl vector
    function [1600:0] proc_path(input [PROC_NUM - 1:0] dl_vec);
        integer index;
        begin
            index = proc_index(dl_vec);
            case (index)
                0 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_46_1_proc_U0";
                end
                1 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_55_2_proc_U0";
                end
                2 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0";
                end
                3 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_1_U0";
                end
                4 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_U0";
                end
                5 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0";
                end
                6 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0";
                end
                7 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_Block_entry1_proc_U0";
                end
                8 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0";
                end
                9 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0";
                end
                10 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0";
                end
                11 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_Block_entry1_proc_U0";
                end
                12 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0";
                end
                13 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0";
                end
                14 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0";
                end
                15 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0";
                end
                16 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0";
                end
                17 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0";
                end
                18 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_U0";
                end
                19 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0";
                end
                20 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0";
                end
                21 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0";
                end
                22 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0";
                end
                23 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7235_proc_U0";
                end
                24 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.ConvertShiftAbs_U0";
                end
                25 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7237_proc_U0";
                end
                26 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.erode_0_0_600_800_0_3_3_1_1_2_2_U0";
                end
                27 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7239_proc_U0";
                end
                28 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.dilate_0_0_600_800_0_3_3_1_1_2_2_U0";
                end
                29 : begin
                    proc_path = "stereolbm_axis_cambm_stereolbm_axis_cambm.xfMat2AXIvideo_8_0_600_800_1_2_U0";
                end
                default : begin
                    proc_path = "unknown";
                end
            endcase
        end
    endfunction

    // print the headlines of deadlock detection
    task print_dl_head;
        begin
            $display("\n//////////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", $time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            fp = $fopen("deadlock_db.dat", "w");
        end
    endtask

    // print the start of a cycle
    task print_cycle_start(input reg [1600:0] proc_path, input integer cycle_id);
        begin
            $display("/////////////////////////");
            $display("// Dependence cycle %0d:", cycle_id);
            $display("// (1): Process: %0s", proc_path);
            $fdisplay(fp, "Dependence_Cycle_ID %0d", cycle_id);
            $fdisplay(fp, "Dependence_Process_ID 1");
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print the end of deadlock detection
    task print_dl_end(input integer num, input integer record_time);
        begin
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// Totally %0d cycles detected!", num);
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", record_time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            $fdisplay(fp, "Dependence_Cycle_Number %0d", num);
            $fclose(fp);
        end
    endtask

    // print one proc component in the cycle
    task print_cycle_proc_comp(input reg [1600:0] proc_path, input integer cycle_comp_id);
        begin
            $display("// (%0d): Process: %0s", cycle_comp_id, proc_path);
            $fdisplay(fp, "Dependence_Process_ID %0d", cycle_comp_id);
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print one channel component in the cycle
    task print_cycle_chan_comp(input [PROC_NUM - 1:0] dl_vec1, input [PROC_NUM - 1:0] dl_vec2);
        reg [1696:0] chan_path;
        integer index1;
        integer index2;
        begin
            index1 = proc_index(dl_vec1);
            index2 = proc_index(dl_vec2);
            case (index1)
                0 : begin
                    case(index2)
                    9: begin
                        if (~irA_r_fix_U.i_full_n & Loop_VITIS_LOOP_46_1_proc_U0.ap_done & ap_done_reg_0 & ~irA_r_fix_U.t_read) begin
                            if (~irA_r_fix_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.irA_r_fix_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.irA_r_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~irA_r_fix_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.irA_r_fix_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.irA_r_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~cameraMA_r_fix_U.i_full_n & Loop_VITIS_LOOP_46_1_proc_U0.ap_done & ap_done_reg_0 & ~cameraMA_r_fix_U.t_read) begin
                            if (~cameraMA_r_fix_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.cameraMA_r_fix_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.cameraMA_r_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~cameraMA_r_fix_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.cameraMA_r_fix_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.cameraMA_r_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    5: begin
                        if (~irA_l_fix_U.i_full_n & Loop_VITIS_LOOP_46_1_proc_U0.ap_done & ap_done_reg_0 & ~irA_l_fix_U.t_read) begin
                            if (~irA_l_fix_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.irA_l_fix_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.irA_l_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~irA_l_fix_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.irA_l_fix_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.irA_l_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~cameraMA_l_fix_U.i_full_n & Loop_VITIS_LOOP_46_1_proc_U0.ap_done & ap_done_reg_0 & ~cameraMA_l_fix_U.t_read) begin
                            if (~cameraMA_l_fix_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.cameraMA_l_fix_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.cameraMA_l_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~cameraMA_l_fix_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.cameraMA_l_fix_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.cameraMA_l_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin
                        if (ap_sync_Loop_VITIS_LOOP_46_1_proc_U0_ap_ready & Loop_VITIS_LOOP_46_1_proc_U0.ap_idle & ~ap_sync_Loop_VITIS_LOOP_55_2_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_55_2_proc_U0'");
                        end
                    end
                    2: begin
                        if (ap_sync_Loop_VITIS_LOOP_46_1_proc_U0_ap_ready & Loop_VITIS_LOOP_46_1_proc_U0.ap_idle & ~ap_sync_Block_for_end72_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                        end
                    end
                    23: begin
                        if (ap_sync_Loop_VITIS_LOOP_46_1_proc_U0_ap_ready & Loop_VITIS_LOOP_46_1_proc_U0.ap_idle & ~ap_sync_Block_for_end7235_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7235_proc_U0'");
                        end
                    end
                    25: begin
                        if (ap_sync_Loop_VITIS_LOOP_46_1_proc_U0_ap_ready & Loop_VITIS_LOOP_46_1_proc_U0.ap_idle & ~ap_sync_Block_for_end7237_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7237_proc_U0'");
                        end
                    end
                    27: begin
                        if (ap_sync_Loop_VITIS_LOOP_46_1_proc_U0_ap_ready & Loop_VITIS_LOOP_46_1_proc_U0.ap_idle & ~ap_sync_Block_for_end7239_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7239_proc_U0'");
                        end
                    end
                    endcase
                end
                1 : begin
                    case(index2)
                    9: begin
                        if (~distC_r_fix_U.i_full_n & Loop_VITIS_LOOP_55_2_proc_U0.ap_done & ap_done_reg_1 & ~distC_r_fix_U.t_read) begin
                            if (~distC_r_fix_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.distC_r_fix_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.distC_r_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~distC_r_fix_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.distC_r_fix_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.distC_r_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    5: begin
                        if (~distC_l_fix_U.i_full_n & Loop_VITIS_LOOP_55_2_proc_U0.ap_done & ap_done_reg_1 & ~distC_l_fix_U.t_read) begin
                            if (~distC_l_fix_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.distC_l_fix_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.distC_l_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~distC_l_fix_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.distC_l_fix_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.distC_l_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (ap_sync_Loop_VITIS_LOOP_55_2_proc_U0_ap_ready & Loop_VITIS_LOOP_55_2_proc_U0.ap_idle & ~ap_sync_Loop_VITIS_LOOP_46_1_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_46_1_proc_U0'");
                        end
                    end
                    2: begin
                        if (ap_sync_Loop_VITIS_LOOP_55_2_proc_U0_ap_ready & Loop_VITIS_LOOP_55_2_proc_U0.ap_idle & ~ap_sync_Block_for_end72_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                        end
                    end
                    23: begin
                        if (ap_sync_Loop_VITIS_LOOP_55_2_proc_U0_ap_ready & Loop_VITIS_LOOP_55_2_proc_U0.ap_idle & ~ap_sync_Block_for_end7235_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7235_proc_U0'");
                        end
                    end
                    25: begin
                        if (ap_sync_Loop_VITIS_LOOP_55_2_proc_U0_ap_ready & Loop_VITIS_LOOP_55_2_proc_U0.ap_idle & ~ap_sync_Block_for_end7237_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7237_proc_U0'");
                        end
                    end
                    27: begin
                        if (ap_sync_Loop_VITIS_LOOP_55_2_proc_U0_ap_ready & Loop_VITIS_LOOP_55_2_proc_U0.ap_idle & ~ap_sync_Block_for_end7239_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7239_proc_U0'");
                        end
                    end
                    endcase
                end
                2 : begin
                    case(index2)
                    0: begin
                        if (ap_sync_Block_for_end72_proc_U0_ap_ready & Block_for_end72_proc_U0.ap_idle & ~ap_sync_Loop_VITIS_LOOP_46_1_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_46_1_proc_U0'");
                        end
                    end
                    1: begin
                        if (ap_sync_Block_for_end72_proc_U0_ap_ready & Block_for_end72_proc_U0.ap_idle & ~ap_sync_Loop_VITIS_LOOP_55_2_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_55_2_proc_U0'");
                        end
                    end
                    23: begin
                        if (ap_sync_Block_for_end72_proc_U0_ap_ready & Block_for_end72_proc_U0.ap_idle & ~ap_sync_Block_for_end7235_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7235_proc_U0'");
                        end
                    end
                    25: begin
                        if (ap_sync_Block_for_end72_proc_U0_ap_ready & Block_for_end72_proc_U0.ap_idle & ~ap_sync_Block_for_end7237_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7237_proc_U0'");
                        end
                    end
                    27: begin
                        if (ap_sync_Block_for_end72_proc_U0_ap_ready & Block_for_end72_proc_U0.ap_idle & ~ap_sync_Block_for_end7239_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7239_proc_U0'");
                        end
                    end
                    endcase
                end
                3 : begin
                    case(index2)
                    2: begin
                        if (~imgL_in_rows_c59_channel_U.if_empty_n & AXIvideo2xfMat_8_0_600_800_1_2_1_U0.ap_idle & ~imgL_in_rows_c59_channel_U.if_write) begin
                            if (~imgL_in_rows_c59_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c59_channel_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c59_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgL_in_rows_c59_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c59_channel_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c59_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~imgL_in_cols_c60_channel_U.if_empty_n & AXIvideo2xfMat_8_0_600_800_1_2_1_U0.ap_idle & ~imgL_in_cols_c60_channel_U.if_write) begin
                            if (~imgL_in_cols_c60_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c60_channel_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c60_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgL_in_cols_c60_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c60_channel_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c60_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    6: begin
                        if (~AXIvideo2xfMat_8_0_600_800_1_2_1_U0.grp_AXIvideo2xfMat_8_0_600_800_1_2_1_Pipeline_loop_col_zxi2mat_fu_205.imgL_in_data_blk_n) begin
                            if (~imgL_in_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgL_in_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AXIvideo2xfMat_8_0_600_800_1_2_1_U0.imgL_in_rows_c_blk_n) begin
                            if (~imgL_in_rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgL_in_rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AXIvideo2xfMat_8_0_600_800_1_2_1_U0.imgL_in_cols_c_blk_n) begin
                            if (~imgL_in_cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgL_in_cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0_U.if_full_n & AXIvideo2xfMat_8_0_600_800_1_2_1_U0.ap_start & ~AXIvideo2xfMat_8_0_600_800_1_2_1_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.start_for_remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0',");
                        end
                    end
                    8: begin
                        if (~AXIvideo2xfMat_8_0_600_800_1_2_1_U0.grp_AXIvideo2xfMat_8_0_600_800_1_2_1_Pipeline_loop_col_zxi2mat_fu_205.imgL_in_data_blk_n) begin
                            if (~imgL_in_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgL_in_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    7: begin
                        if (~AXIvideo2xfMat_8_0_600_800_1_2_1_U0.imgL_in_rows_c_blk_n) begin
                            if (~imgL_in_rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_Block_entry1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgL_in_rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_Block_entry1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AXIvideo2xfMat_8_0_600_800_1_2_1_U0.imgL_in_cols_c_blk_n) begin
                            if (~imgL_in_cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_Block_entry1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgL_in_cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_Block_entry1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                4 : begin
                    case(index2)
                    2: begin
                        if (~imgR_in_rows_c61_channel_U.if_empty_n & AXIvideo2xfMat_8_0_600_800_1_2_U0.ap_idle & ~imgR_in_rows_c61_channel_U.if_write) begin
                            if (~imgR_in_rows_c61_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c61_channel_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c61_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgR_in_rows_c61_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c61_channel_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c61_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~imgR_in_cols_c62_channel_U.if_empty_n & AXIvideo2xfMat_8_0_600_800_1_2_U0.ap_idle & ~imgR_in_cols_c62_channel_U.if_write) begin
                            if (~imgR_in_cols_c62_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c62_channel_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c62_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgR_in_cols_c62_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c62_channel_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c62_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    10: begin
                        if (~AXIvideo2xfMat_8_0_600_800_1_2_U0.grp_AXIvideo2xfMat_8_0_600_800_1_2_Pipeline_loop_col_zxi2mat_fu_205.imgR_in_data_blk_n) begin
                            if (~imgR_in_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgR_in_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AXIvideo2xfMat_8_0_600_800_1_2_U0.imgR_in_rows_c_blk_n) begin
                            if (~imgR_in_rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgR_in_rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AXIvideo2xfMat_8_0_600_800_1_2_U0.imgR_in_cols_c_blk_n) begin
                            if (~imgR_in_cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgR_in_cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0_U.if_full_n & AXIvideo2xfMat_8_0_600_800_1_2_U0.ap_start & ~AXIvideo2xfMat_8_0_600_800_1_2_U0.real_start & (trans_in_cnt_1 == trans_out_cnt_1) & ~start_for_remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.start_for_remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0',");
                        end
                    end
                    12: begin
                        if (~AXIvideo2xfMat_8_0_600_800_1_2_U0.grp_AXIvideo2xfMat_8_0_600_800_1_2_Pipeline_loop_col_zxi2mat_fu_205.imgR_in_data_blk_n) begin
                            if (~imgR_in_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgR_in_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    11: begin
                        if (~AXIvideo2xfMat_8_0_600_800_1_2_U0.imgR_in_rows_c_blk_n) begin
                            if (~imgR_in_rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_Block_entry1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgR_in_rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_Block_entry1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AXIvideo2xfMat_8_0_600_800_1_2_U0.imgR_in_cols_c_blk_n) begin
                            if (~imgR_in_cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_Block_entry1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgR_in_cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_Block_entry1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                5 : begin
                    case(index2)
                    0: begin
                        if (~cameraMA_l_fix_U.t_empty_n & InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0.ap_idle & ~cameraMA_l_fix_U.i_write) begin
                            if (~cameraMA_l_fix_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.cameraMA_l_fix_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_46_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.cameraMA_l_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~cameraMA_l_fix_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.cameraMA_l_fix_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_46_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.cameraMA_l_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~irA_l_fix_U.t_empty_n & InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0.ap_idle & ~irA_l_fix_U.i_write) begin
                            if (~irA_l_fix_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.irA_l_fix_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_46_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.irA_l_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~irA_l_fix_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.irA_l_fix_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_46_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.irA_l_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin
                        if (~distC_l_fix_U.t_empty_n & InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0.ap_idle & ~distC_l_fix_U.i_write) begin
                            if (~distC_l_fix_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.distC_l_fix_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_55_2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.distC_l_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~distC_l_fix_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.distC_l_fix_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_55_2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.distC_l_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    2: begin
                        if (~mapxLMat_rows_U.if_empty_n & InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0.ap_idle & ~mapxLMat_rows_U.if_write) begin
                            if (~mapxLMat_rows_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_rows_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_rows_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapxLMat_rows_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_rows_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_rows_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~mapxLMat_cols_U.if_empty_n & InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0.ap_idle & ~mapxLMat_cols_U.if_write) begin
                            if (~mapxLMat_cols_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_cols_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_cols_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapxLMat_cols_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_cols_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_cols_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    6: begin
                        if (~InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0.grp_xFInitUndistortRectifyMapInverseKernel_fu_40.grp_xFInitUndistortRectifyMapInverseKernel_Pipeline_loop_height_loop_width_fu_152.mapxRMat_data_blk_n) begin
                            if (~mapxLMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapxLMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0.grp_xFInitUndistortRectifyMapInverseKernel_fu_40.grp_xFInitUndistortRectifyMapInverseKernel_Pipeline_loop_height_loop_width_fu_152.mapyRMat_data_blk_n) begin
                            if (~mapyLMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapyLMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapyLMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapyLMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapyLMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapyLMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    8: begin
                        if (~InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0.grp_xFInitUndistortRectifyMapInverseKernel_fu_40.grp_xFInitUndistortRectifyMapInverseKernel_Pipeline_loop_height_loop_width_fu_152.mapxRMat_data_blk_n) begin
                            if (~mapxLMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapxLMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0.grp_xFInitUndistortRectifyMapInverseKernel_fu_40.grp_xFInitUndistortRectifyMapInverseKernel_Pipeline_loop_height_loop_width_fu_152.mapyRMat_data_blk_n) begin
                            if (~mapyLMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapyLMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapyLMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapyLMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapyLMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapyLMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                6 : begin
                    case(index2)
                    3: begin
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_Block_entry1_proc_U0.p_src_mat_rows_blk_n) begin
                            if (~imgL_in_rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgL_in_rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_Block_entry1_proc_U0.p_src_mat_cols_blk_n) begin
                            if (~imgL_in_cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgL_in_cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_Pipeline_loop_width_fu_104.imgL_in_data_blk_n) begin
                            if (~imgL_in_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgL_in_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0_U.if_empty_n & remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.ap_idle & ~start_for_remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.start_for_remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_1_U0',");
                        end
                    end
                    13: begin
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_Pipeline_loop_width_fu_104.leftRemappedMat_data_blk_n) begin
                            if (~leftRemappedMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~leftRemappedMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    5: begin
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_Pipeline_loop_width_fu_104.mapxLMat_data_blk_n) begin
                            if (~mapxLMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapxLMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_Pipeline_loop_width_fu_104.mapyLMat_data_blk_n) begin
                            if (~mapyLMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapyLMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapyLMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapyLMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapyLMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapyLMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                7 : begin
                    case(index2)
                    3: begin
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_Block_entry1_proc_U0.p_src_mat_rows_blk_n) begin
                            if (~imgL_in_rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgL_in_rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_Block_entry1_proc_U0.p_src_mat_cols_blk_n) begin
                            if (~imgL_in_cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgL_in_cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                8 : begin
                    case(index2)
                    3: begin
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_Pipeline_loop_width_fu_104.imgL_in_data_blk_n) begin
                            if (~imgL_in_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgL_in_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgL_in_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    13: begin
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_Pipeline_loop_width_fu_104.leftRemappedMat_data_blk_n) begin
                            if (~leftRemappedMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~leftRemappedMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    5: begin
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_Pipeline_loop_width_fu_104.mapxLMat_data_blk_n) begin
                            if (~mapxLMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapxLMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxLMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_Pipeline_loop_width_fu_104.mapyLMat_data_blk_n) begin
                            if (~mapyLMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapyLMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapyLMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapyLMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapyLMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapyLMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    7: begin
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.rows_loc_channel_U.if_empty_n & remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0.ap_idle & ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.rows_loc_channel_U.if_write) begin
                            if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.rows_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.rows_loc_channel_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_Block_entry1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.rows_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.rows_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.rows_loc_channel_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_Block_entry1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.rows_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.cols_loc_channel_U.if_empty_n & remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0.ap_idle & ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.cols_loc_channel_U.if_write) begin
                            if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.cols_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.cols_loc_channel_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_Block_entry1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.cols_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.cols_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.cols_loc_channel_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_Block_entry1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.cols_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                9 : begin
                    case(index2)
                    0: begin
                        if (~cameraMA_r_fix_U.t_empty_n & InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0.ap_idle & ~cameraMA_r_fix_U.i_write) begin
                            if (~cameraMA_r_fix_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.cameraMA_r_fix_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_46_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.cameraMA_r_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~cameraMA_r_fix_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.cameraMA_r_fix_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_46_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.cameraMA_r_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~irA_r_fix_U.t_empty_n & InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0.ap_idle & ~irA_r_fix_U.i_write) begin
                            if (~irA_r_fix_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.irA_r_fix_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_46_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.irA_r_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~irA_r_fix_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.irA_r_fix_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_46_1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.irA_r_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin
                        if (~distC_r_fix_U.t_empty_n & InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0.ap_idle & ~distC_r_fix_U.i_write) begin
                            if (~distC_r_fix_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.distC_r_fix_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_55_2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.distC_r_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~distC_r_fix_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'stereolbm_axis_cambm_stereolbm_axis_cambm.distC_r_fix_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_55_2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.distC_r_fix_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    2: begin
                        if (~mapxRMat_rows_U.if_empty_n & InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0.ap_idle & ~mapxRMat_rows_U.if_write) begin
                            if (~mapxRMat_rows_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_rows_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_rows_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapxRMat_rows_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_rows_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_rows_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~mapxRMat_cols_U.if_empty_n & InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0.ap_idle & ~mapxRMat_cols_U.if_write) begin
                            if (~mapxRMat_cols_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_cols_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_cols_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapxRMat_cols_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_cols_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_cols_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    10: begin
                        if (~InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0.grp_xFInitUndistortRectifyMapInverseKernel_fu_40.grp_xFInitUndistortRectifyMapInverseKernel_Pipeline_loop_height_loop_width_fu_152.mapxRMat_data_blk_n) begin
                            if (~mapxRMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapxRMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0.grp_xFInitUndistortRectifyMapInverseKernel_fu_40.grp_xFInitUndistortRectifyMapInverseKernel_Pipeline_loop_height_loop_width_fu_152.mapyRMat_data_blk_n) begin
                            if (~mapyRMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapyRMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapyRMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapyRMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapyRMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapyRMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    12: begin
                        if (~InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0.grp_xFInitUndistortRectifyMapInverseKernel_fu_40.grp_xFInitUndistortRectifyMapInverseKernel_Pipeline_loop_height_loop_width_fu_152.mapxRMat_data_blk_n) begin
                            if (~mapxRMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapxRMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0.grp_xFInitUndistortRectifyMapInverseKernel_fu_40.grp_xFInitUndistortRectifyMapInverseKernel_Pipeline_loop_height_loop_width_fu_152.mapyRMat_data_blk_n) begin
                            if (~mapyRMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapyRMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapyRMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapyRMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapyRMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapyRMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                10 : begin
                    case(index2)
                    4: begin
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_Block_entry1_proc_U0.p_src_mat_rows_blk_n) begin
                            if (~imgR_in_rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgR_in_rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_Block_entry1_proc_U0.p_src_mat_cols_blk_n) begin
                            if (~imgR_in_cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgR_in_cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_Pipeline_loop_width_fu_104.imgR_in_data_blk_n) begin
                            if (~imgR_in_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgR_in_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0_U.if_empty_n & remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.ap_idle & ~start_for_remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.start_for_remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_U0',");
                        end
                    end
                    13: begin
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_Pipeline_loop_width_fu_104.rightRemappedMat_data_blk_n) begin
                            if (~rightRemappedMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rightRemappedMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    9: begin
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_Pipeline_loop_width_fu_104.mapxRMat_data_blk_n) begin
                            if (~mapxRMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapxRMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_Pipeline_loop_width_fu_104.mapyRMat_data_blk_n) begin
                            if (~mapyRMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapyRMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapyRMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapyRMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapyRMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapyRMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                11 : begin
                    case(index2)
                    4: begin
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_Block_entry1_proc_U0.p_src_mat_rows_blk_n) begin
                            if (~imgR_in_rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgR_in_rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_Block_entry1_proc_U0.p_src_mat_cols_blk_n) begin
                            if (~imgR_in_cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgR_in_cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                12 : begin
                    case(index2)
                    4: begin
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_Pipeline_loop_width_fu_104.imgR_in_data_blk_n) begin
                            if (~imgR_in_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgR_in_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.AXIvideo2xfMat_8_0_600_800_1_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.imgR_in_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    13: begin
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_Pipeline_loop_width_fu_104.rightRemappedMat_data_blk_n) begin
                            if (~rightRemappedMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rightRemappedMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    9: begin
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_Pipeline_loop_width_fu_104.mapxRMat_data_blk_n) begin
                            if (~mapxRMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapxRMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapxRMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0.grp_xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_Pipeline_loop_width_fu_104.mapyRMat_data_blk_n) begin
                            if (~mapyRMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapyRMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapyRMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~mapyRMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.mapyRMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.InitUndistortRectifyMapInverse_9_5_7_600_800_1_2_2_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.mapyRMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    11: begin
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.rows_loc_channel_U.if_empty_n & remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0.ap_idle & ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.rows_loc_channel_U.if_write) begin
                            if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.rows_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.rows_loc_channel_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_Block_entry1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.rows_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.rows_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.rows_loc_channel_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_Block_entry1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.rows_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.cols_loc_channel_U.if_empty_n & remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0.ap_idle & ~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.cols_loc_channel_U.if_write) begin
                            if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.cols_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.cols_loc_channel_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_Block_entry1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.cols_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.cols_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.cols_loc_channel_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_Block_entry1_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.cols_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                13 : begin
                    case(index2)
                    2: begin
                        if (~leftRemappedMat_rows_U.if_empty_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.ap_idle & ~leftRemappedMat_rows_U.if_write) begin
                            if (~leftRemappedMat_rows_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_rows_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_rows_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~leftRemappedMat_rows_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_rows_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_rows_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~leftRemappedMat_cols_U.if_empty_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.ap_idle & ~leftRemappedMat_cols_U.if_write) begin
                            if (~leftRemappedMat_cols_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_cols_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_cols_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~leftRemappedMat_cols_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_cols_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_cols_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~rightRemappedMat_rows_U.if_empty_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.ap_idle & ~rightRemappedMat_rows_U.if_write) begin
                            if (~rightRemappedMat_rows_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_rows_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_rows_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rightRemappedMat_rows_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_rows_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_rows_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~rightRemappedMat_cols_U.if_empty_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.ap_idle & ~rightRemappedMat_cols_U.if_write) begin
                            if (~rightRemappedMat_cols_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_cols_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_cols_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rightRemappedMat_cols_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_cols_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_cols_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~bmState_preFilterCap_U.if_empty_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.ap_idle & ~bmState_preFilterCap_U.if_write) begin
                            if (~bmState_preFilterCap_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.bmState_preFilterCap_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.bmState_preFilterCap_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bmState_preFilterCap_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.bmState_preFilterCap_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.bmState_preFilterCap_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~bmState_textureThreshold_U.if_empty_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.ap_idle & ~bmState_textureThreshold_U.if_write) begin
                            if (~bmState_textureThreshold_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.bmState_textureThreshold_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.bmState_textureThreshold_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bmState_textureThreshold_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.bmState_textureThreshold_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.bmState_textureThreshold_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~bmState_uniquenessRatio_U.if_empty_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.ap_idle & ~bmState_uniquenessRatio_U.if_write) begin
                            if (~bmState_uniquenessRatio_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.bmState_uniquenessRatio_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.bmState_uniquenessRatio_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bmState_uniquenessRatio_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.bmState_uniquenessRatio_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.bmState_uniquenessRatio_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    6: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0.grp_xFSobelFilter3x3_0_3_600_800_1_0_4_1_2_2_2_1_6_800_false_s_fu_36.grp_xFSobelFilter3x3_Pipeline_Clear_Row_Loop_fu_148.rightRemappedMat_data_blk_n) begin
                            if (~leftRemappedMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~leftRemappedMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    8: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0.grp_xFSobelFilter3x3_0_3_600_800_1_0_4_1_2_2_2_1_6_800_false_s_fu_36.grp_xFSobelFilter3x3_Pipeline_Clear_Row_Loop_fu_148.rightRemappedMat_data_blk_n) begin
                            if (~leftRemappedMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~leftRemappedMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.leftRemappedMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    10: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_U0.grp_xFSobelFilter3x3_0_3_600_800_1_0_4_1_2_2_2_1_6_800_false_s_fu_36.grp_xFSobelFilter3x3_Pipeline_Clear_Row_Loop_fu_148.rightRemappedMat_data_blk_n) begin
                            if (~rightRemappedMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rightRemappedMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    12: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_U0.grp_xFSobelFilter3x3_0_3_600_800_1_0_4_1_2_2_2_1_6_800_false_s_fu_36.grp_xFSobelFilter3x3_Pipeline_Clear_Row_Loop_fu_148.rightRemappedMat_data_blk_n) begin
                            if (~rightRemappedMat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rightRemappedMat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.remap_128_1_0_7_0_600_800_1_false_2_2_2_2_U0.xFRemapLI_0_0_1_7_128_600_800_1_2_2_2_2_false_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.rightRemappedMat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    24: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0.grp_xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_Pipeline_VITIS_LOOP_fu_46.img_disp16u_data_blk_n) begin
                            if (~img_disp16u_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp16u_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.ConvertShiftAbs_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp16u_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_disp16u_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp16u_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.ConvertShiftAbs_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp16u_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_ConvertShiftAbs_U0_U.if_full_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.ap_start & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.real_start & (trans_in_cnt_4 == trans_out_cnt_4) & ~start_for_ConvertShiftAbs_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.start_for_ConvertShiftAbs_U0_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.ConvertShiftAbs_U0',");
                        end
                    end
                    endcase
                end
                14 : begin
                    case(index2)
                    19: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.sbmstate_preFilterCap_c18_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c18_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c18_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.height_c22_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c22_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c22_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.width_c27_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c27_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c27_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFImageClip_600_800_1_2_4_0_3_0_800_U0_U.if_full_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.ap_start & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.real_start & (trans_in_cnt_2 == trans_out_cnt_2) & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFImageClip_600_800_1_2_4_0_3_0_800_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFImageClip_600_800_1_2_4_0_3_0_800_U0_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0',");
                        end
                    end
                    16: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.sbmstate_preFilterCap_c19_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c19_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c19_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.height_c24_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c24_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c24_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.width_c29_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c29_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c29_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFImageClip_600_800_1_2_4_0_3_0_800_4_U0_U.if_full_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.ap_start & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.real_start & (trans_in_cnt_2 == trans_out_cnt_2) & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFImageClip_600_800_1_2_4_0_3_0_800_4_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFImageClip_600_800_1_2_4_0_3_0_800_4_U0_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0',");
                        end
                    end
                    21: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.sbmstate_textureThreshold_c_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_textureThreshold_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_textureThreshold_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_textureThreshold_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_textureThreshold_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_textureThreshold_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_textureThreshold_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.sbmstate_uniquenessRatio_c_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_uniquenessRatio_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_uniquenessRatio_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_uniquenessRatio_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_uniquenessRatio_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_uniquenessRatio_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_uniquenessRatio_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFSADBlockMatching_U0_U.if_full_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.ap_start & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.real_start & (trans_in_cnt_2 == trans_out_cnt_2) & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFSADBlockMatching_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFSADBlockMatching_U0_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0',");
                        end
                    end
                    20: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.height_c21_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c21_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c21_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.width_c26_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c26_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c26_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFReadOutStream_600_800_1_2_4_0_3_800_U0_U.if_full_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.ap_start & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.real_start & (trans_in_cnt_2 == trans_out_cnt_2) & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFReadOutStream_600_800_1_2_4_0_3_800_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFReadOutStream_600_800_1_2_4_0_3_800_U0_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0',");
                        end
                    end
                    17: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.height_c23_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c23_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c23_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.width_c28_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c28_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c28_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFReadOutStream_600_800_1_2_4_0_3_800_5_U0_U.if_full_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.ap_start & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.real_start & (trans_in_cnt_2 == trans_out_cnt_2) & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFReadOutStream_600_800_1_2_4_0_3_800_5_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFReadOutStream_600_800_1_2_4_0_3_800_5_U0_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0',");
                        end
                    end
                    15: begin
                        if (StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.ap_sync_entry_proc_U0_ap_ready & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.ap_idle & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.ap_sync_Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0'");
                        end
                    end
                    18: begin
                        if (StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.ap_sync_entry_proc_U0_ap_ready & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0.ap_idle & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.ap_sync_Sobel_0_3_0_3_600_800_1_false_2_2_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_U0'");
                        end
                    end
                    endcase
                end
                15 : begin
                    case(index2)
                    16: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0.grp_xFSobelFilter3x3_0_3_600_800_1_0_4_1_2_2_2_1_6_800_false_s_fu_36.grp_xFSobelFilter3x3_Pipeline_Col_Loop_fu_157.in_sobel_x_i_data_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    17: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0.grp_xFSobelFilter3x3_0_3_600_800_1_0_4_1_2_2_2_1_6_800_false_s_fu_36.grp_xFSobelFilter3x3_Pipeline_Col_Loop_fu_157.in_sobel_y_i_data_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    14: begin
                        if (StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.ap_sync_Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0_ap_ready & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0.ap_idle & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                        end
                    end
                    18: begin
                        if (StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.ap_sync_Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0_ap_ready & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0.ap_idle & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.ap_sync_Sobel_0_3_0_3_600_800_1_false_2_2_2_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_U0'");
                        end
                    end
                    endcase
                end
                16 : begin
                    case(index2)
                    15: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0.grp_xFImageClip_600_800_1_2_4_0_3_0_800_4_Pipeline_loop_col_clip_fu_108.in_sobel_x_data_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    21: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0.grp_xFImageClip_600_800_1_2_4_0_3_0_800_4_Pipeline_loop_col_clip_fu_108.left_clipped_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.left_clipped_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.left_clipped_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.left_clipped_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.left_clipped_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.left_clipped_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.left_clipped_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0.sbmstate_preFilterCap_c_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0.height_c20_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c20_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c20_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0.width_c25_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c25_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c25_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    14: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0.sbmstate_preFilterCap_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c19_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c19_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0.height_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c24_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c24_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c24_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c24_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0.width_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c29_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c29_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c29_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c29_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFImageClip_600_800_1_2_4_0_3_0_800_4_U0_U.if_empty_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0.ap_idle & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFImageClip_600_800_1_2_4_0_3_0_800_4_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFImageClip_600_800_1_2_4_0_3_0_800_4_U0_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0',");
                        end
                    end
                    endcase
                end
                17 : begin
                    case(index2)
                    15: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0.grp_xFReadOutStream_600_800_1_2_4_0_3_800_5_Pipeline_loop_col_clip_fu_62.in_sobel_y_i4_data_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    14: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0.height_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c23_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c23_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c23_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c23_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0.width_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c28_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c28_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c28_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c28_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFReadOutStream_600_800_1_2_4_0_3_800_5_U0_U.if_empty_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0.ap_idle & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFReadOutStream_600_800_1_2_4_0_3_800_5_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFReadOutStream_600_800_1_2_4_0_3_800_5_U0_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0',");
                        end
                    end
                    20: begin
                        if (ap_done_reg_12 & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0.ap_done & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_12 & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0.ap_done & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0'");
                        end
                    end
                    endcase
                end
                18 : begin
                    case(index2)
                    19: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_U0.grp_xFSobelFilter3x3_0_3_600_800_1_0_4_1_2_2_2_1_6_800_false_s_fu_36.grp_xFSobelFilter3x3_Pipeline_Col_Loop_fu_157.in_sobel_x_i_data_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_1_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_1_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    20: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_U0.grp_xFSobelFilter3x3_0_3_600_800_1_0_4_1_2_2_2_1_6_800_false_s_fu_36.grp_xFSobelFilter3x3_Pipeline_Col_Loop_fu_157.in_sobel_y_i_data_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_1_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_1_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    14: begin
                        if (StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.ap_sync_Sobel_0_3_0_3_600_800_1_false_2_2_2_U0_ap_ready & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_U0.ap_idle & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.ap_sync_entry_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                        end
                    end
                    15: begin
                        if (StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.ap_sync_Sobel_0_3_0_3_600_800_1_false_2_2_2_U0_ap_ready & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_U0.ap_idle & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.ap_sync_Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_3_U0'");
                        end
                    end
                    endcase
                end
                19 : begin
                    case(index2)
                    18: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0.grp_xFImageClip_600_800_1_2_4_0_3_0_800_Pipeline_loop_col_clip_fu_74.in_sobel_x_data_1_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_1_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_1_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_x_data_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    21: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0.grp_xFImageClip_600_800_1_2_4_0_3_0_800_Pipeline_loop_col_clip_fu_74.right_clipped_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.right_clipped_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.right_clipped_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.right_clipped_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.right_clipped_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.right_clipped_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.right_clipped_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    14: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0.sbmstate_preFilterCap_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c18_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c18_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0.height_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c22_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c22_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c22_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c22_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0.width_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c27_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c27_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c27_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c27_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFImageClip_600_800_1_2_4_0_3_0_800_U0_U.if_empty_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0.ap_idle & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFImageClip_600_800_1_2_4_0_3_0_800_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFImageClip_600_800_1_2_4_0_3_0_800_U0_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0',");
                        end
                    end
                    endcase
                end
                20 : begin
                    case(index2)
                    18: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0.grp_xFReadOutStream_600_800_1_2_4_0_3_800_Pipeline_loop_col_clip_fu_62.in_sobel_y_i_data_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_1_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_1_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.Sobel_0_3_0_3_600_800_1_false_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.in_sobel_y_data_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    14: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0.height_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c21_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c21_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c21_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c21_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0.width_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c26_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c26_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c26_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c26_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFReadOutStream_600_800_1_2_4_0_3_800_U0_U.if_empty_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0.ap_idle & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFReadOutStream_600_800_1_2_4_0_3_800_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFReadOutStream_600_800_1_2_4_0_3_800_U0_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0',");
                        end
                    end
                    17: begin
                        if (ap_done_reg_13 & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0.ap_done & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_13 & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0.ap_done & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0'");
                        end
                    end
                    endcase
                end
                21 : begin
                    case(index2)
                    16: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0.grp_xFSADBlockMatching_Pipeline_loop_row_loop_mux_loop_col_fu_106.left_clipped_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.left_clipped_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.left_clipped_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.left_clipped_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.left_clipped_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.left_clipped_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.left_clipped_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0.state_preFilterCap_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_preFilterCap_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0.height_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c20_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c20_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c20_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c20_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0.width_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c25_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c25_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c25_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c25_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_4_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0.grp_xFSADBlockMatching_Pipeline_loop_row_loop_mux_loop_col_fu_106.right_clipped_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.right_clipped_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.right_clipped_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.right_clipped_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.right_clipped_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.right_clipped_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFImageClip_600_800_1_2_4_0_3_0_800_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.right_clipped_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    22: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0.grp_xFSADBlockMatching_Pipeline_loop_row_loop_mux_loop_col_fu_106.p_disp_strm_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.p_disp_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.p_disp_strm_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.p_disp_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.p_disp_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.p_disp_strm_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.p_disp_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0.height_c_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0.width_c_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0_U.if_full_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0.ap_start & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0.real_start & (trans_in_cnt_3 == trans_out_cnt_3) & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0',");
                        end
                    end
                    14: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0.state_textureThreshold_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_textureThreshold_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_textureThreshold_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_textureThreshold_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_textureThreshold_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_textureThreshold_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_textureThreshold_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0.state_uniquenessRatio_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_uniquenessRatio_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_uniquenessRatio_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_uniquenessRatio_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_uniquenessRatio_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_uniquenessRatio_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.sbmstate_uniquenessRatio_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFSADBlockMatching_U0_U.if_empty_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0.ap_idle & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFSADBlockMatching_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFSADBlockMatching_U0_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.entry_proc_U0',");
                        end
                    end
                    endcase
                end
                22 : begin
                    case(index2)
                    21: begin
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0.width_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0.height_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.height_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0.grp_xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_Pipeline_VITIS_LOOP_fu_46.p_disp_strm_blk_n) begin
                            if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.p_disp_strm_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.p_disp_strm_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.p_disp_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.p_disp_strm_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.p_disp_strm_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.p_disp_strm_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0_U.if_empty_n & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0.ap_idle & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.start_for_xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFSADBlockMatching_U0',");
                        end
                    end
                    17: begin
                        if (ap_done_reg_14 & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0.ap_done & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_5_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_14 & StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFFindStereoCorrespondenceLBMNO_Loop_VITIS_LOOP_816_1_proc13_U0.ap_done & ~StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0.grp_xFFindStereoCorrespondenceLBMNO_fu_76.xFReadOutStream_600_800_1_2_4_0_3_800_U0'");
                        end
                    end
                    endcase
                end
                23 : begin
                    case(index2)
                    0: begin
                        if (ap_sync_Block_for_end7235_proc_U0_ap_ready & Block_for_end7235_proc_U0.ap_idle & ~ap_sync_Loop_VITIS_LOOP_46_1_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_46_1_proc_U0'");
                        end
                    end
                    1: begin
                        if (ap_sync_Block_for_end7235_proc_U0_ap_ready & Block_for_end7235_proc_U0.ap_idle & ~ap_sync_Loop_VITIS_LOOP_55_2_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_55_2_proc_U0'");
                        end
                    end
                    2: begin
                        if (ap_sync_Block_for_end7235_proc_U0_ap_ready & Block_for_end7235_proc_U0.ap_idle & ~ap_sync_Block_for_end72_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                        end
                    end
                    25: begin
                        if (ap_sync_Block_for_end7235_proc_U0_ap_ready & Block_for_end7235_proc_U0.ap_idle & ~ap_sync_Block_for_end7237_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7237_proc_U0'");
                        end
                    end
                    27: begin
                        if (ap_sync_Block_for_end7235_proc_U0_ap_ready & Block_for_end7235_proc_U0.ap_idle & ~ap_sync_Block_for_end7239_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7239_proc_U0'");
                        end
                    end
                    endcase
                end
                24 : begin
                    case(index2)
                    13: begin
                        if (~ConvertShiftAbs_U0.grp_ConvertShiftAbs_Pipeline_loop_width_fu_38.img_disp16u_data_blk_n) begin
                            if (~img_disp16u_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp16u_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp16u_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_disp16u_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp16u_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp16u_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_ConvertShiftAbs_U0_U.if_empty_n & ConvertShiftAbs_U0.ap_idle & ~start_for_ConvertShiftAbs_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.start_for_ConvertShiftAbs_U0_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.StereoBM_15_128_16_0_2_600_800_1_false_2_2_2_U0',");
                        end
                    end
                    26: begin
                        if (~ConvertShiftAbs_U0.grp_ConvertShiftAbs_Pipeline_loop_width_fu_38.img_disp8u_data_blk_n) begin
                            if (~img_disp8u_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.erode_0_0_600_800_0_3_3_1_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_disp8u_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.erode_0_0_600_800_0_3_3_1_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                25 : begin
                    case(index2)
                    0: begin
                        if (ap_sync_Block_for_end7237_proc_U0_ap_ready & Block_for_end7237_proc_U0.ap_idle & ~ap_sync_Loop_VITIS_LOOP_46_1_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_46_1_proc_U0'");
                        end
                    end
                    1: begin
                        if (ap_sync_Block_for_end7237_proc_U0_ap_ready & Block_for_end7237_proc_U0.ap_idle & ~ap_sync_Loop_VITIS_LOOP_55_2_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_55_2_proc_U0'");
                        end
                    end
                    2: begin
                        if (ap_sync_Block_for_end7237_proc_U0_ap_ready & Block_for_end7237_proc_U0.ap_idle & ~ap_sync_Block_for_end72_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                        end
                    end
                    23: begin
                        if (ap_sync_Block_for_end7237_proc_U0_ap_ready & Block_for_end7237_proc_U0.ap_idle & ~ap_sync_Block_for_end7235_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7235_proc_U0'");
                        end
                    end
                    27: begin
                        if (ap_sync_Block_for_end7237_proc_U0_ap_ready & Block_for_end7237_proc_U0.ap_idle & ~ap_sync_Block_for_end7239_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7239_proc_U0'");
                        end
                    end
                    endcase
                end
                26 : begin
                    case(index2)
                    23: begin
                        if (~img_disp8u_rows_U.if_empty_n & erode_0_0_600_800_0_3_3_1_1_2_2_U0.ap_idle & ~img_disp8u_rows_U.if_write) begin
                            if (~img_disp8u_rows_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_rows_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7235_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_rows_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_disp8u_rows_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_rows_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7235_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_rows_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~img_disp8u_cols_U.if_empty_n & erode_0_0_600_800_0_3_3_1_1_2_2_U0.ap_idle & ~img_disp8u_cols_U.if_write) begin
                            if (~img_disp8u_cols_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_cols_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7235_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_cols_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_disp8u_cols_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_cols_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7235_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_cols_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    24: begin
                        if (~erode_0_0_600_800_0_3_3_1_1_2_2_U0.grp_xferode_600_800_1_0_1_2_2_0_801_3_3_s_fu_34.grp_xferode_600_800_1_0_1_2_2_0_801_3_3_Pipeline_Col_Loop_fu_155.img_disp8u_data_blk_n) begin
                            if (~img_disp8u_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.ConvertShiftAbs_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_disp8u_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.ConvertShiftAbs_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    28: begin
                        if (~erode_0_0_600_800_0_3_3_1_1_2_2_U0.grp_xferode_600_800_1_0_1_2_2_0_801_3_3_s_fu_34.grp_xferode_600_800_1_0_1_2_2_0_801_3_3_Pipeline_Col_Loop_fu_155.img_disp8u_erode_data_blk_n) begin
                            if (~img_disp8u_erode_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_erode_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.dilate_0_0_600_800_0_3_3_1_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_erode_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_disp8u_erode_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_erode_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.dilate_0_0_600_800_0_3_3_1_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_erode_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                27 : begin
                    case(index2)
                    0: begin
                        if (ap_sync_Block_for_end7239_proc_U0_ap_ready & Block_for_end7239_proc_U0.ap_idle & ~ap_sync_Loop_VITIS_LOOP_46_1_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_46_1_proc_U0'");
                        end
                    end
                    1: begin
                        if (ap_sync_Block_for_end7239_proc_U0_ap_ready & Block_for_end7239_proc_U0.ap_idle & ~ap_sync_Loop_VITIS_LOOP_55_2_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Loop_VITIS_LOOP_55_2_proc_U0'");
                        end
                    end
                    2: begin
                        if (ap_sync_Block_for_end7239_proc_U0_ap_ready & Block_for_end7239_proc_U0.ap_idle & ~ap_sync_Block_for_end72_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end72_proc_U0'");
                        end
                    end
                    23: begin
                        if (ap_sync_Block_for_end7239_proc_U0_ap_ready & Block_for_end7239_proc_U0.ap_idle & ~ap_sync_Block_for_end7235_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7235_proc_U0'");
                        end
                    end
                    25: begin
                        if (ap_sync_Block_for_end7239_proc_U0_ap_ready & Block_for_end7239_proc_U0.ap_idle & ~ap_sync_Block_for_end7237_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7237_proc_U0'");
                        end
                    end
                    endcase
                end
                28 : begin
                    case(index2)
                    25: begin
                        if (~img_disp8u_erode_rows_U.if_empty_n & dilate_0_0_600_800_0_3_3_1_1_2_2_U0.ap_idle & ~img_disp8u_erode_rows_U.if_write) begin
                            if (~img_disp8u_erode_rows_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_erode_rows_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7237_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_erode_rows_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_disp8u_erode_rows_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_erode_rows_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7237_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_erode_rows_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~img_disp8u_erode_cols_U.if_empty_n & dilate_0_0_600_800_0_3_3_1_1_2_2_U0.ap_idle & ~img_disp8u_erode_cols_U.if_write) begin
                            if (~img_disp8u_erode_cols_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_erode_cols_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7237_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_erode_cols_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_disp8u_erode_cols_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_erode_cols_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7237_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_erode_cols_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    26: begin
                        if (~dilate_0_0_600_800_0_3_3_1_1_2_2_U0.grp_xfdilate_600_800_1_0_1_2_2_0_801_3_3_s_fu_34.grp_xfdilate_600_800_1_0_1_2_2_0_801_3_3_Pipeline_Col_Loop_fu_155.img_disp8u_erode_data_blk_n) begin
                            if (~img_disp8u_erode_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_erode_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.erode_0_0_600_800_0_3_3_1_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_erode_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_disp8u_erode_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_erode_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.erode_0_0_600_800_0_3_3_1_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_erode_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    29: begin
                        if (~dilate_0_0_600_800_0_3_3_1_1_2_2_U0.grp_xfdilate_600_800_1_0_1_2_2_0_801_3_3_s_fu_34.grp_xfdilate_600_800_1_0_1_2_2_0_801_3_3_Pipeline_Col_Loop_fu_155.img_disp8u_dilate_data_blk_n) begin
                            if (~img_disp8u_dilate_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_dilate_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.xfMat2AXIvideo_8_0_600_800_1_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_dilate_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_disp8u_dilate_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_dilate_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.xfMat2AXIvideo_8_0_600_800_1_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_dilate_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                29 : begin
                    case(index2)
                    27: begin
                        if (~img_disp8u_dilate_rows_U.if_empty_n & xfMat2AXIvideo_8_0_600_800_1_2_U0.ap_idle & ~img_disp8u_dilate_rows_U.if_write) begin
                            if (~img_disp8u_dilate_rows_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_dilate_rows_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7239_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_dilate_rows_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_disp8u_dilate_rows_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_dilate_rows_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7239_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_dilate_rows_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~img_disp8u_dilate_cols_U.if_empty_n & xfMat2AXIvideo_8_0_600_800_1_2_U0.ap_idle & ~img_disp8u_dilate_cols_U.if_write) begin
                            if (~img_disp8u_dilate_cols_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_dilate_cols_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7239_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_dilate_cols_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_disp8u_dilate_cols_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_dilate_cols_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.Block_for_end7239_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_dilate_cols_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    28: begin
                        if (~xfMat2AXIvideo_8_0_600_800_1_2_U0.grp_xfMat2AXIvideo_8_0_600_800_1_2_Pipeline_loop_col_mat2axi_fu_86.img_disp8u_dilate_data_blk_n) begin
                            if (~img_disp8u_dilate_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_dilate_data_U' written by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.dilate_0_0_600_800_0_3_3_1_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_dilate_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_disp8u_dilate_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_dilate_data_U' read by process 'stereolbm_axis_cambm_stereolbm_axis_cambm.dilate_0_0_600_800_0_3_3_1_1_2_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path stereolbm_axis_cambm_stereolbm_axis_cambm.img_disp8u_dilate_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
            endcase
        end
    endtask

    // report
    initial begin : report_deadlock
        integer cycle_id;
        integer cycle_comp_id;
        integer record_time;
        wait (dl_reset == 1);
        cycle_id = 1;
        record_time = 0;
        while (1) begin
            @ (negedge dl_clock);
            case (CS_fsm)
                ST_DL_DETECTED: begin
                    cycle_comp_id = 2;
                    if (dl_detect_reg != dl_done_reg) begin
                        if (dl_done_reg == 'b0) begin
                            print_dl_head;
                            record_time = $time;
                        end
                        print_cycle_start(proc_path(origin), cycle_id);
                        cycle_id = cycle_id + 1;
                    end
                    else begin
                        print_dl_end((cycle_id - 1),record_time);
                        @(negedge dl_clock);
                        @(negedge dl_clock);
                        $finish;
                    end
                end
                ST_DL_REPORT: begin
                    if ((|(dl_in_vec)) & ~(|(dl_in_vec & origin_reg))) begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                        print_cycle_proc_comp(proc_path(dl_in_vec), cycle_comp_id);
                        cycle_comp_id = cycle_comp_id + 1;
                    end
                    else begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                    end
                end
            endcase
        end
    end
 
